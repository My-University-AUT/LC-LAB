`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//  
// Made by: Ali Nowrouzi and Ahmad Foroughi 
// 
// Create Date:    17:23:14 11/01/2020 
//////////////////////////////////////////////////////////////////////////////////
module X_NOR_2(input A,B,C, output out
    );
	xnor(out,A,B,C);
endmodule
